`ifndef C_ROUNDING_TRANSACTION
`define C_ROUNDING_TRANSACTION

class c_rounding_transaction;
int	y_rounding;
int cb_rounding;
int cr_rounding;
endclass : c_rounding_transaction

`endif
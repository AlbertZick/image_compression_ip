`ifndef C_SEQUENCER
`define C_SEQUENCER

typedef uvm_sequencer #(c_random_item) c_sequencer;

`endif
# vsim -novopt -c "+num_sequence=1000" top -do "run -all;exit;" -l log.svh 
# Start time: 11:19:35 on Aug 29,2018
# ** Warning: (vsim-8891) All optimizations are turned off because the -novopt switch is in effect. This will cause your simulation to run very slowly. If you are using this switch to preserve visibility for Debug or PLI features please see the User's Manual section on Preserving Object Visibility with vopt.
# 
# //  Questa Sim
# //  Version 10.4e win32 Apr  9 2016
# //
# //  Copyright 1991-2016 Mentor Graphics Corporation
# //  All Rights Reserved.
# //
# //  THIS WORK CONTAINS TRADE SECRET AND PROPRIETARY INFORMATION
# //  WHICH IS THE PROPERTY OF MENTOR GRAPHICS CORPORATION OR ITS
# //  LICENSORS AND IS SUBJECT TO LICENSE TERMS.
# //  THIS DOCUMENT CONTAINS TRADE SECRETS AND COMMERCIAL OR FINANCIAL
# //  INFORMATION THAT ARE PRIVILEGED, CONFIDENTIAL, AND EXEMPT FROM
# //  DISCLOSURE UNDER THE FREEDOM OF INFORMATION ACT, 5 U.S.C. SECTION 552.
# //  FURTHERMORE, THIS INFORMATION IS PROHIBITED FROM DISCLOSURE UNDER
# //  THE TRADE SECRETS ACT, 18 U.S.C. SECTION 1905.
# //
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.top
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.pkg_uvm_test
# Loading sv_std.std
# Loading mtiUvm.uvm_pkg
# Loading work.pkg_uvm_test
# Loading work.top
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.if_dut
# Loading work.if_dut
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_dut
# Loading work.m_dut
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_small_ip
# Loading work.m_small_ip
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.convert_int_into_float
# Loading work.convert_int_into_float
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.abs_25_bits
# Loading work.abs_25_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.mux_2_1
# Loading work.mux_2_1
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.cong_25bits
# Loading work.cong_25bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.full_adder
# Loading work.full_adder
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_1_25bits
# Loading work.shift_left_1_25bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.adder_unsign_8_bits
# Loading work.adder_unsign_8_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_nadd_9_sign_bits
# Loading work.sub_nadd_9_sign_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.convert_color_space_Y
# Loading work.convert_color_space_Y
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.FP
# Loading work.FP
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.small_ALU
# Loading work.small_ALU
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.exponent_difference
# Loading work.exponent_difference
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_right
# Loading work.shift_right
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.big_ALU
# Loading work.big_ALU
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.demux_1_4
# Loading work.demux_1_4
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.demux_1_2
# Loading work.demux_1_2
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_nadd_25_sign_bits
# Loading work.sub_nadd_25_sign_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_24x24_bits
# Loading work.multiplier_24x24_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_12x12_bits
# Loading work.multiplier_12x12_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_6x6_bits
# Loading work.multiplier_6x6_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.add_24_bits
# Loading work.add_24_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.add_48_bits
# Loading work.add_48_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.divider_24x24_bits
# Loading work.divider_24x24_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.mux_4_1
# Loading work.mux_4_1
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.abs
# Loading work.abs
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_nadd_49_sign_bits
# Loading work.sub_nadd_49_sign_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.inc_or_dec
# Loading work.inc_or_dec
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_or_right
# Loading work.shift_left_or_right
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_24_bits
# Loading work.shift_left_24_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_12_bits
# Loading work.shift_left_12_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_6_bits
# Loading work.shift_left_6_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.shift_left_1_bit
# Loading work.shift_left_1_bit
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.adder_unsign_6_bits
# Loading work.adder_unsign_6_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_unsign_6_bits
# Loading work.sub_unsign_6_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.FP_control
# Loading work.FP_control
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.rounding
# Loading work.rounding
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.convert_color_space_Cb
# Loading work.convert_color_space_Cb
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.convert_color_space_Cr
# Loading work.convert_color_space_Cr
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.control_convertion
# Loading work.control_convertion
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.mem_YCbCr
# Loading work.mem_YCbCr
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.convert_float_into_int
# Loading work.convert_float_into_int
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.adjust_significand
# Loading work.adjust_significand
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.decide_on_rounding
# Loading work.decide_on_rounding
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.control_DCT
# Loading work.control_DCT
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.dct_2_D
# Loading work.dct_2_D
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.dct
# Loading work.dct
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_2
# Loading work.multiplier_2
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.dich_trai_1
# Loading work.dich_trai_1
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_6
# Loading work.multiplier_6
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_8
# Loading work.multiplier_8
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_14
# Loading work.multiplier_14
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.tru_25bits
# Loading work.tru_25bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_15
# Loading work.multiplier_15
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_16
# Loading work.multiplier_16
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_19
# Loading work.multiplier_19
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_30
# Loading work.multiplier_30
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_35
# Loading work.multiplier_35
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_36
# Loading work.multiplier_36
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.multiplier_39
# Loading work.multiplier_39
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.dieu_chinh
# Loading work.dieu_chinh
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.mem_8x8
# Loading work.mem_8x8
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.counter_8_state
# Loading work.counter_8_state
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.D_flipflop
# Loading work.D_flipflop
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.delay_1_clk
# Loading work.delay_1_clk
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.control_quatization
# Loading work.control_quatization
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.Y_quantization
# Loading work.Y_quantization
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.Chrominance_quantization
# Loading work.Chrominance_quantization
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_control_encoder
# Loading work.m_control_encoder
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_luminance_component_encoder
# Loading work.m_luminance_component_encoder
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_bin_counter
# Loading work.m_bin_counter
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.FF
# Loading work.FF
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.mem_64
# Loading work.mem_64
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_zigzac_table
# Loading work.m_zigzac_table
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_delay_28_clock
# Loading work.m_delay_28_clock
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_ZZk_comparator
# Loading work.m_ZZk_comparator
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_K_comparator
# Loading work.m_K_comparator
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_reg_R
# Loading work.m_reg_R
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_R_comparator
# Loading work.m_R_comparator
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_encode_luminance_ac
# Loading work.m_encode_luminance_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_calc_ac_addl_bits
# Loading work.m_calc_ac_addl_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_calc_ac_category
# Loading work.m_calc_ac_category
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_nadd_11_sign_bits
# Loading work.sub_nadd_11_sign_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_luminance_huff_code_ac
# Loading work.m_luminance_huff_code_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_luminance_ext_hm_code_ac
# Loading work.m_luminance_ext_hm_code_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.adder_unsign_5_bits
# Loading work.adder_unsign_5_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_encode_luminance_dc
# Loading work.m_encode_luminance_dc
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_dc_diff
# Loading work.m_dc_diff
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_calc_dc_category
# Loading work.m_calc_dc_category
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.sub_nadd_12_sign_bits
# Loading work.sub_nadd_12_sign_bits
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_luminance_huff_code_dc
# Loading work.m_luminance_huff_code_dc
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_luminance_ext_hm_code_dc
# Loading work.m_luminance_ext_hm_code_dc
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_control_v2
# Loading work.m_control_v2
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_chrominance_component_encoder
# Loading work.m_chrominance_component_encoder
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_encode_chrominance_ac
# Loading work.m_encode_chrominance_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_chrominance_huff_code_ac
# Loading work.m_chrominance_huff_code_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_chrominance_ext_hm_code_ac
# Loading work.m_chrominance_ext_hm_code_ac
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_encode_chrominance_dc
# Loading work.m_encode_chrominance_dc
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_chrominance_huff_code_dc
# Loading work.m_chrominance_huff_code_dc
# Refreshing F:/MyProjects/TruongTran/AMCC/UVM_projects/Image_compression/uvm_test_v2/work.m_chrominance_ext_hm_code_dc
# Loading work.m_chrominance_ext_hm_code_dc
# Loading mtiUvm.questa_uvm_pkg
# Loading F:/MyPrograms/questasim_10.4e/uvm-1.1d\win32\uvm_dpi.dll
# run -all
# ----------------------------------------------------------------
# UVM-1.1d
# (C) 2007-2013 Mentor Graphics Corporation
# (C) 2007-2013 Cadence Design Systems, Inc.
# (C) 2006-2013 Synopsys, Inc.
# (C) 2011-2013 Cypress Semiconductor Corp.
# ----------------------------------------------------------------
# 
#   ***********       IMPORTANT RELEASE NOTES         ************
# 
#   You are using a version of the UVM library that has been compiled
#   with `UVM_NO_DEPRECATED undefined.
#   See http://www.eda.org/svdb/view.php?id=3313 for more details.
# 
#   You are using a version of the UVM library that has been compiled
#   with `UVM_OBJECT_MUST_HAVE_CONSTRUCTOR undefined.
#   See http://www.eda.org/svdb/view.php?id=3770 for more details.
# 
#       (Specify +UVM_NO_RELNOTES to turn off this notice)
# 
# UVM_INFO verilog_src/questa_uvm_pkg-1.2/src/questa_uvm_pkg.sv(215) @ 0: reporter [Questa UVM] QUESTA_UVM-1.2.3
# UVM_INFO verilog_src/questa_uvm_pkg-1.2/src/questa_uvm_pkg.sv(217) @ 0: reporter [Questa UVM]  questa_uvm::init(+struct)
# UVM_INFO @ 0: reporter [RNTST] Running test c_random_test...
# UVM_INFO c_scoreboard.svh(251) @ 8000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 8000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 8000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(251) @ 15680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 15680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 15680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 17960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 17960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 17960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 17960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 17960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 17960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 17960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 17960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 17960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 21400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 21400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 21400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 23360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 23360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 23360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 25640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 25640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 25640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 25640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 25640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 25640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 25640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 25640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 25640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 29080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 29080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 29080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 31040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 31040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 31040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 33320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 33320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 33320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 33320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 33320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 33320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 33320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 33320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 33320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 36760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 36760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 36760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 38720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 38720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 38720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 41000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 41000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 41000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 41000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 41000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 41000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 41000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 41000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 41000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 44440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 44440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 44440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 46400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 46400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 46400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 48680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 48680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 48680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 48680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 48680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 48680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 48680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 48680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 48680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 52120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 52120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 52120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 54080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 54080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 54080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 56360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 56360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 56360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 56360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 56360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 56360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 56360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 56360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 56360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 59800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 59800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 59800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 61760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 61760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 61760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 64040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 64040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 64040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 64040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 64040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 64040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 64040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 64040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 64040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 67480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 67480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 67480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 69440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 69440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 69440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 71720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 71720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 71720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 71720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 71720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 71720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 71720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 71720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 71720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 75160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 75160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 75160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 77120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 77120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 77120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 79400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 79400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 79400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 79400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 79400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 79400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 79400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 79400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 79400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 82840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 82840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 82840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 84800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 84800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 84800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 87080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 87080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 87080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 87080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 87080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 87080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 87080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 87080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 87080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 90520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 90520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 90520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 92480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 92480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 92480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 94760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 94760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 94760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 94760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 94760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 94760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 94760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 94760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 94760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 98200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 98200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 98200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 100160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 100160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 100160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 102440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 102440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 102440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 102440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 102440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 102440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 102440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 102440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 102440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 105880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 105880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 105880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 107840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 107840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 107840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 110120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 110120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 110120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 110120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 110120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 110120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 110120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 110120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 110120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 113560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 113560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 113560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 115520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 115520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 115520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 117800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 117800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 117800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 117800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 117800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 117800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 117800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 117800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 117800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 121240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 121240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 121240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 123200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 123200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 123200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 125480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 125480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 125480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 125480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 125480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 125480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 125480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 125480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 125480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 128920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 128920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 128920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 130880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 130880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 130880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 133160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 133160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 133160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 133160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 133160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 133160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 133160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 133160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 133160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 136600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 136600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 136600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 138560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 138560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 138560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 140840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 140840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 140840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 140840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 140840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 140840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 140840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 140840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 140840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 144280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 144280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 144280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 146240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 146240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 146240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 148520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 148520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 148520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 148520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 148520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 148520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 148520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 148520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 148520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 151960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 151960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 151960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 153920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 153920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 153920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 156200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 156200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 156200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 156200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 156200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 156200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 156200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 156200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 156200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 159640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 159640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 159640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 161600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 161600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 161600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 163880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 163880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 163880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 163880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 163880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 163880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 163880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 163880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 163880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 167320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 167320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 167320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 169280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 169280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 169280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 171560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 171560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 171560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 171560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 171560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 171560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 171560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 171560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 171560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 175000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 175000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 175000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 176960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 176960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 176960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 179240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 179240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 179240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 179240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 179240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 179240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 179240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 179240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 179240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 182680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 182680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 182680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 184640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 184640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 184640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 186920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 186920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 186920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 186920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 186920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 186920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 186920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 186920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 186920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 190360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 190360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 190360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 192320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 192320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 192320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 194600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 194600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 194600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 194600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 194600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 194600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 194600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 194600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 194600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 198040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 198040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 198040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 200000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 200000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 200000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 202280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 202280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 202280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 202280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 202280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 202280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 202280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 202280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 202280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 205720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 205720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 205720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 207680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 207680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 207680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 209960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 209960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 209960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 209960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 209960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 209960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 209960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 209960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 209960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 213400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 213400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 213400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 215360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 215360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 215360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 217640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 217640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 217640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 217640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 217640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 217640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 217640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 217640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 217640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 221080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 221080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 221080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 223040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 223040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 223040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 225320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 225320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 225320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 225320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 225320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 225320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 225320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 225320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 225320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 228760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 228760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 228760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 230720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 230720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 230720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 233000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 233000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 233000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 233000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 233000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 233000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 233000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 233000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 233000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 236440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 236440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 236440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 238400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 238400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 238400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 240680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 240680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 240680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 240680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 240680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 240680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 240680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 240680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 240680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 244120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 244120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 244120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 246080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 246080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 246080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 248360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 248360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 248360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 248360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 248360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 248360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 248360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 248360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 248360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 251800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 251800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 251800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 253760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 253760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 253760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 256040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 256040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 256040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 256040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 256040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 256040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 256040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 256040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 256040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 259480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 259480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 259480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 261440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 261440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 261440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 263720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 263720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 263720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 263720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 263720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 263720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 263720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 263720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 263720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 267160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 267160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 267160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 269120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 269120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 269120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 271400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 271400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 271400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 271400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 271400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 271400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 271400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 271400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 271400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 274840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 274840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 274840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 276800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 276800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 276800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 279080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 279080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 279080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 279080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 279080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 279080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 279080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 279080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 279080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 282520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 282520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 282520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 284480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 284480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 284480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 286760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 286760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 286760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 286760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 286760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 286760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 286760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 286760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 286760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 290200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 290200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 290200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 292160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 292160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 292160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 294440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 294440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 294440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 294440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 294440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 294440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 294440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 294440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 294440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 297880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 297880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 297880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 299840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 299840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 299840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 302120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 302120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 302120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 302120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 302120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 302120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 302120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 302120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 302120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 305560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 305560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 305560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 307520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 307520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 307520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 309800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 309800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 309800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 309800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 309800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 309800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 309800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 309800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 309800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 313240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 313240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 313240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 315200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 315200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 315200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 317480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 317480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 317480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 317480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 317480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 317480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 317480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 317480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 317480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 320920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 320920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 320920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 322880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 322880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 322880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 325160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 325160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 325160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 325160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 325160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 325160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 325160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 325160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 325160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 328600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 328600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 328600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 330560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 330560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 330560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 332840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 332840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 332840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 332840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 332840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 332840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 332840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 332840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 332840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 336280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 336280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 336280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 338240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 338240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 338240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 340520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 340520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 340520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 340520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 340520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 340520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 340520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 340520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 340520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 343960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 343960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 343960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 345920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 345920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 345920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 348200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 348200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 348200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 348200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 348200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 348200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 348200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 348200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 348200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 351640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 351640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 351640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 353600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 353600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 353600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 355880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 355880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 355880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 355880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 355880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 355880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 355880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 355880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 355880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 359320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 359320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 359320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 361280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 361280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 361280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 363560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 363560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 363560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 363560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 363560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 363560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 363560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 363560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 363560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 367000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 367000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 367000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 368960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 368960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 368960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 371240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 371240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 371240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 371240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 371240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 371240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 371240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 371240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 371240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 374680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 374680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 374680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 376640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 376640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 376640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 378920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 378920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 378920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 378920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 378920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 378920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 378920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 378920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 378920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 382360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 382360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 382360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 384320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 384320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 384320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 386600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 386600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 386600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 386600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 386600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 386600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 386600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 386600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 386600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 390040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 390040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 390040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 392000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 392000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 392000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 394280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 394280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 394280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 394280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 394280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 394280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 394280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 394280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 394280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 397720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 397720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 397720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 399680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 399680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 399680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 401960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 401960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 401960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 401960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 401960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 401960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 401960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 401960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 401960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 405400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 405400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 405400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 407360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 407360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 407360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 409640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 409640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 409640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 409640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 409640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 409640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 409640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 409640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 409640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 413080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 413080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 413080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 415040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 415040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 415040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 417320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 417320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 417320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 417320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 417320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 417320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 417320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 417320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 417320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 420760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 420760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 420760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 422720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 422720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 422720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 425000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 425000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 425000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 425000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 425000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 425000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 425000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 425000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 425000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 428440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 428440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 428440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 430400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 430400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 430400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 432680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 432680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 432680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 432680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 432680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 432680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 432680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 432680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 432680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 436120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 436120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 436120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 438080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 438080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 438080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 440360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 440360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 440360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 440360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 440360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 440360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 440360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 440360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 440360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 443800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 443800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 443800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 445760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 445760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 445760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 448040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 448040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 448040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 448040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 448040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 448040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 448040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 448040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 448040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 451480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 451480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 451480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 453440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 453440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 453440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 455720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 455720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 455720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 455720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 455720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 455720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 455720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 455720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 455720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 459160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 459160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 459160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 461120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 461120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 461120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 463400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 463400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 463400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 463400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 463400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 463400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 463400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 463400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 463400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 466840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 466840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 466840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 468800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 468800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 468800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 471080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 471080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 471080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 471080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 471080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 471080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 471080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 471080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 471080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 474520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 474520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 474520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 476480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 476480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 476480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 478760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 478760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 478760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 478760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 478760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 478760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 478760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 478760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 478760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 482200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 482200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 482200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 484160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 484160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 484160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 486440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 486440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 486440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 486440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 486440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 486440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 486440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 486440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 486440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 489880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 489880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 489880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 491840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 491840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 491840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 494120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 494120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 494120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 494120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 494120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 494120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 494120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 494120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 494120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 497560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 497560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 497560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 499520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 499520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 499520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 501800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 501800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 501800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 501800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 501800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 501800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 501800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 501800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 501800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 505240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 505240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 505240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 507200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 507200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 507200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 509480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 509480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 509480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 509480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 509480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 509480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 509480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 509480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 509480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 512920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 512920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 512920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 514880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 514880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 514880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 517160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 517160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 517160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 517160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 517160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 517160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 517160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 517160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 517160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 520600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 520600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 520600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 522560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 522560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 522560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 524840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 524840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 524840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 524840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 524840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 524840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 524840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 524840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 524840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 528280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 528280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 528280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 530240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 530240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 530240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 532520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 532520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 532520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 532520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 532520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 532520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 532520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 532520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 532520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 535960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 535960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 535960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 537920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 537920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 537920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 540200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 540200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 540200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 540200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 540200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 540200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 540200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 540200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 540200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 543640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 543640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 543640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 545600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 545600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 545600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 547880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 547880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 547880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 547880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 547880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 547880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 547880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 547880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 547880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 551320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 551320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 551320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 553280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 553280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 553280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 555560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 555560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 555560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 555560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 555560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 555560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 555560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 555560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 555560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 559000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 559000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 559000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 560960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 560960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 560960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 563240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 563240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 563240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 563240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 563240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 563240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 563240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 563240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 563240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 566680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 566680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 566680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 568640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 568640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 568640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 570920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 570920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 570920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 570920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 570920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 570920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 570920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 570920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 570920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 574360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 574360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 574360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 576320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 576320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 576320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 578600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 578600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 578600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 578600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 578600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 578600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 578600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 578600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 578600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 582040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 582040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 582040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 584000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 584000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 584000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 586280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 586280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 586280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 586280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 586280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 586280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 586280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 586280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 586280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 589720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 589720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 589720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 591680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 591680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 591680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 593960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 593960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 593960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 593960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 593960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 593960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 593960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 593960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 593960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 597400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 597400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 597400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 599360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 599360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 599360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 601640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 601640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 601640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 601640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 601640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 601640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 601640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 601640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 601640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 605080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 605080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 605080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 607040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 607040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 607040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 609320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 609320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 609320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 609320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 609320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 609320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 609320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 609320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 609320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 612760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 612760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 612760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 614720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 614720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 614720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 617000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 617000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 617000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 617000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 617000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 617000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 617000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 617000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 617000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 620440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 620440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 620440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 622400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 622400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 622400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 624680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 624680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 624680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 624680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 624680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 624680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 624680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 624680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 624680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 628120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 628120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 628120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 630080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 630080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 630080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 632360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 632360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 632360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 632360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 632360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 632360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 632360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 632360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 632360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 635800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 635800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 635800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 637760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 637760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 637760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 640040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 640040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 640040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 640040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 640040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 640040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 640040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 640040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 640040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 643480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 643480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 643480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 645440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 645440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 645440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 647720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 647720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 647720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 647720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 647720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 647720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 647720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 647720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 647720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 651160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 651160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 651160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 653120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 653120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 653120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 655400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 655400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 655400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 655400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 655400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 655400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 655400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 655400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 655400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 658840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 658840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 658840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 660800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 660800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 660800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 663080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 663080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 663080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 663080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 663080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 663080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 663080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 663080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 663080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 666520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 666520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 666520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 668480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 668480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 668480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 670760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 670760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 670760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 670760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 670760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 670760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 670760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 670760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 670760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 674200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 674200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 674200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 676160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 676160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 676160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 678440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 678440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 678440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 678440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 678440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 678440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 678440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 678440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 678440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 681880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 681880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 681880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 683840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 683840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 683840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 686120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 686120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 686120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 686120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 686120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 686120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 686120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 686120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 686120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 689560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 689560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 689560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 691520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 691520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 691520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 693800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 693800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 693800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 693800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 693800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 693800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 693800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 693800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 693800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 697240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 697240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 697240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 699200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 699200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 699200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 701480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 701480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 701480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 701480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 701480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 701480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 701480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 701480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 701480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 704920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 704920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 704920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 706880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 706880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 706880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 709160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 709160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 709160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 709160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 709160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 709160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 709160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 709160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 709160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 712600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 712600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 712600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 714560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 714560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 714560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 716840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 716840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 716840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 716840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 716840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 716840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 716840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 716840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 716840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 720280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 720280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 720280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 722240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 722240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 722240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 724520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 724520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 724520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 724520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 724520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 724520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 724520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 724520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 724520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 727960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 727960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 727960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 729920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 729920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 729920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 732200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 732200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 732200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 732200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 732200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 732200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 732200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 732200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 732200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 735640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 735640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 735640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 737600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 737600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 737600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 739880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 739880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 739880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 739880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 739880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 739880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 739880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 739880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 739880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 743320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 743320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 743320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 745280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 745280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 745280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 747560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 747560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 747560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 747560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 747560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 747560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 747560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 747560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 747560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 751000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 751000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 751000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 752960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 752960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 752960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 755240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 755240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 755240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 755240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 755240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 755240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 755240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 755240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 755240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 758680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 758680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 758680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 760640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 760640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 760640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 762920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 762920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 762920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 762920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 762920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 762920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 762920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 762920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 762920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 766360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 766360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 766360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 768320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 768320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 768320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 770600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 770600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 770600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 770600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 770600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 770600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 770600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 770600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 770600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 774040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 774040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 774040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 776000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 776000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 776000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 778280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 778280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 778280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 778280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 778280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 778280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 778280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 778280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 778280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 781720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 781720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 781720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 783680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 783680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 783680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 785960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 785960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 785960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 785960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 785960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 785960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 785960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 785960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 785960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 789400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 789400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 789400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 791360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 791360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 791360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 793640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 793640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 793640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 793640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 793640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 793640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 793640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 793640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 793640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 797080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 797080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 797080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 799040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 799040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 799040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 801320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 801320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 801320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 801320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 801320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 801320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 801320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 801320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 801320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 804760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 804760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 804760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 806720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 806720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 806720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 809000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 809000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 809000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 809000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 809000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 809000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 809000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 809000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 809000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 812440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 812440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 812440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 814400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 814400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 814400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 816680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 816680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 816680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 816680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 816680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 816680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 816680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 816680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 816680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 820120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 820120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 820120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 822080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 822080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 822080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 824360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 824360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 824360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 824360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 824360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 824360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 824360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 824360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 824360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 827800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 827800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 827800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 829760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 829760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 829760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 832040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 832040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 832040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 832040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 832040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 832040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 832040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 832040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 832040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 835480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 835480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 835480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 837440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 837440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 837440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 839720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 839720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 839720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 839720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 839720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 839720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 839720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 839720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 839720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 843160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 843160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 843160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 845120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 845120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 845120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 847400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 847400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 847400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 847400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 847400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 847400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 847400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 847400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 847400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 850840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 850840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 850840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 852800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 852800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 852800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 855080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 855080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 855080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 855080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 855080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 855080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 855080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 855080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 855080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 858520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 858520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 858520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 860480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 860480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 860480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 862760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 862760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 862760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 862760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 862760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 862760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 862760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 862760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 862760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 866200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 866200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 866200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 868160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 868160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 868160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 870440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 870440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 870440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 870440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 870440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 870440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 870440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 870440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 870440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 873880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 873880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 873880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 875840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 875840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 875840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 878120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 878120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 878120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 878120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 878120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 878120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 878120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 878120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 878120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 881560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 881560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 881560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 883520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 883520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 883520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 885800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 885800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 885800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 885800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 885800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 885800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 885800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 885800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 885800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 889240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 889240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 889240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 891200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 891200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 891200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 893480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 893480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 893480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 893480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 893480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 893480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 893480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 893480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 893480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 896920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 896920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 896920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 898880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 898880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 898880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 901160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 901160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 901160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 901160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 901160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 901160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 901160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 901160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 901160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 904600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 904600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 904600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 906560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 906560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 906560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 908840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 908840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 908840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 908840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 908840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 908840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 908840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 908840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 908840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 912280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 912280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 912280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 914240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 914240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 914240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 916520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 916520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 916520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 916520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 916520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 916520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 916520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 916520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 916520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 919960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 919960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 919960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 921920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 921920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 921920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 924200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 924200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 924200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 924200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 924200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 924200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 924200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 924200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 924200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 927640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 927640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 927640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 929600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 929600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 929600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 931880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 931880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 931880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 931880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 931880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 931880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 931880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 931880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 931880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 935320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 935320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 935320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 937280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 937280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 937280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 939560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 939560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 939560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 939560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 939560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 939560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 939560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 939560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 939560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 943000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 943000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 943000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 944960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 944960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 944960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 947240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 947240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 947240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 947240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 947240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 947240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 947240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 947240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 947240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 950680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 950680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 950680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 952640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 952640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 952640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 954920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 954920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 954920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 954920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 954920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 954920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 954920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 954920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 954920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 958360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 958360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 958360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 960320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 960320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 960320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 962600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 962600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 962600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 962600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 962600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 962600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 962600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 962600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 962600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 966040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 966040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 966040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 968000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 968000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 968000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 970280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 970280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 970280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 970280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 970280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 970280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 970280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 970280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 970280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 973720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 973720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 973720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 975680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 975680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 975680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 977960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 977960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 977960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 977960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 977960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 977960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 977960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 977960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 977960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 981400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 981400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 981400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 983360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 983360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 983360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 985640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 985640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 985640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 985640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 985640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 985640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 985640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 985640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 985640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 989080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 989080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 989080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 991040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 991040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 991040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 993320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 993320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 993320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 993320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 993320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 993320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 993320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 993320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 993320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 996760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 996760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 996760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 998720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 998720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 998720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1001000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1001000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1001000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1001000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1001000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1001000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1001000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1001000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1001000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1004440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1004440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1004440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1006400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1006400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1006400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1008680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1008680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1008680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1008680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1008680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1008680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1008680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1008680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1008680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1012120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1012120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1012120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1014080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1014080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1014080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1016360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1016360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1016360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1016360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1016360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1016360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1016360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1016360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1016360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1019800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1019800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1019800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1021760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1021760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1021760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1024040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1024040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1024040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1024040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1024040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1024040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1024040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1024040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1024040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1027480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1027480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1027480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1029440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1029440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1029440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1031720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1031720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1031720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1031720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1031720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1031720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1031720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1031720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1031720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1035160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1035160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1035160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1037120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1037120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1037120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1039400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1039400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1039400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1039400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1039400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1039400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1039400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1039400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1039400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1042840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1042840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1042840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1044800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1044800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1044800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1047080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1047080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1047080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1047080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1047080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1047080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1047080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1047080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1047080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1050520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1050520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1050520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1052480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1052480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1052480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1054760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1054760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1054760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1054760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1054760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1054760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1054760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1054760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1054760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1058200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1058200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1058200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1060160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1060160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1060160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1062440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1062440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1062440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1062440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1062440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1062440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1062440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1062440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1062440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1065880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1065880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1065880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1067840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1067840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1067840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1070120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1070120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1070120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1070120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1070120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1070120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1070120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1070120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1070120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1073560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1073560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1073560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1075520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1075520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1075520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1077800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1077800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1077800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1077800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1077800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1077800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1077800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1077800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1077800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1081240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1081240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1081240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1083200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1083200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1083200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1085480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1085480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1085480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1085480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1085480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1085480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1085480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1085480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1085480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1088920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1088920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1088920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1090880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1090880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1090880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1093160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1093160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1093160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1093160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1093160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1093160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1093160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1093160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1093160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1096600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1096600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1096600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1098560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1098560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1098560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1100840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1100840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1100840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1100840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1100840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1100840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1100840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1100840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1100840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1104280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1104280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1104280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1106240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1106240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1106240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1108520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1108520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1108520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1108520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1108520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1108520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1108520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1108520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1108520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1111960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1111960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1111960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1113920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1113920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1113920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1116200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1116200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1116200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1116200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1116200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1116200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1116200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1116200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1116200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1119640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1119640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1119640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1121600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1121600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1121600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1123880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1123880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1123880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1123880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1123880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1123880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1123880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1123880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1123880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1127320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1127320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1127320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1129280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1129280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1129280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1131560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1131560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1131560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1131560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1131560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1131560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1131560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1131560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1131560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1135000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1135000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1135000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1136960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1136960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1136960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1139240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1139240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1139240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1139240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1139240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1139240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1139240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1139240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1139240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1142680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1142680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1142680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1144640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1144640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1144640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1146920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1146920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1146920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1146920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1146920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1146920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1146920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1146920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1146920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1150360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1150360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1150360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1152320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1152320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1152320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1154600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1154600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1154600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1154600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1154600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1154600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1154600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1154600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1154600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1158040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1158040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1158040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1160000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1160000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1160000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1162280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1162280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1162280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1162280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1162280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1162280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1162280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1162280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1162280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1165720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1165720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1165720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1167680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1167680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1167680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1169960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1169960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1169960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1169960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1169960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1169960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1169960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1169960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1169960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1173400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1173400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1173400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1175360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1175360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1175360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1177640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1177640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1177640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1177640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1177640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1177640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1177640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1177640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1177640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1181080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1181080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1181080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1183040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1183040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1183040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1185320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1185320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1185320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1185320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1185320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1185320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1185320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1185320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1185320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1188760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1188760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1188760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1190720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1190720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1190720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1193000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1193000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1193000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1193000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1193000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1193000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1193000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1193000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1193000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1196440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1196440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1196440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1198400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1198400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1198400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1200680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1200680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1200680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1200680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1200680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1200680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1200680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1200680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1200680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1204120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1204120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1204120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1206080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1206080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1206080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1208360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1208360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1208360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1208360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1208360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1208360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1208360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1208360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1208360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1211800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1211800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1211800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1213760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1213760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1213760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1216040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1216040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1216040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1216040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1216040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1216040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1216040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1216040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1216040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1219480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1219480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1219480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1221440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1221440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1221440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1223720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1223720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1223720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1223720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1223720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1223720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1223720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1223720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1223720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1227160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1227160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1227160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1229120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1229120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1229120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1231400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1231400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1231400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1231400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1231400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1231400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1231400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1231400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1231400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1234840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1234840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1234840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1236800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1236800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1236800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1239080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1239080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1239080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1239080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1239080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1239080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1239080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1239080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1239080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1242520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1242520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1242520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1244480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1244480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1244480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1246760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1246760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1246760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1246760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1246760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1246760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1246760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1246760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1246760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1250200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1250200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1250200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1252160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1252160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1252160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1254440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1254440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1254440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1254440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1254440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1254440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1254440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1254440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1254440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1257880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1257880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1257880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1259840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1259840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1259840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1262120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1262120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1262120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1262120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1262120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1262120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1262120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1262120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1262120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1265560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1265560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1265560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1267520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1267520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1267520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1269800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1269800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1269800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1269800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1269800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1269800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1269800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1269800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1269800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1273240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1273240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1273240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1275200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1275200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1275200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1277480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1277480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1277480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1277480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1277480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1277480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1277480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1277480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1277480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1280920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1280920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1280920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1282880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1282880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1282880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1285160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1285160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1285160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1285160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1285160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1285160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1285160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1285160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1285160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1288600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1288600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1288600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1290560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1290560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1290560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1292840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1292840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1292840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1292840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1292840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1292840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1292840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1292840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1292840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1296280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1296280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1296280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1298240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1298240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1298240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1300520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1300520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1300520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1300520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1300520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1300520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1300520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1300520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1300520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1303960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1303960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1303960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1305920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1305920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1305920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1308200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1308200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1308200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1308200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1308200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1308200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1308200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1308200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1308200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1311640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1311640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1311640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1313600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1313600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1313600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1315880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1315880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1315880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1315880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1315880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1315880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1315880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1315880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1315880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1319320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1319320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1319320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1321280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1321280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1321280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1323560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1323560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1323560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1323560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1323560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1323560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1323560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1323560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1323560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1327000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1327000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1327000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1328960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1328960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1328960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1331240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1331240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1331240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1331240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1331240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1331240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1331240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1331240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1331240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1334680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1334680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1334680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1336640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1336640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1336640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1338920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1338920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1338920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1338920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1338920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1338920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1338920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1338920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1338920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1342360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1342360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1342360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1344320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1344320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1344320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1346600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1346600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1346600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1346600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1346600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1346600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1346600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1346600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1346600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1350040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1350040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1350040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1352000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1352000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1352000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1354280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1354280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1354280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1354280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1354280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1354280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1354280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1354280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1354280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1357720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1357720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1357720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1359680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1359680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1359680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1361960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1361960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1361960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1361960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1361960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1361960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1361960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1361960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1361960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1365400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1365400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1365400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1367360: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1367360: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1367360: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1369640: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1369640: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1369640: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1369640: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1369640: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1369640: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1369640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1369640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1369640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1373080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1373080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1373080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1375040: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1375040: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1375040: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1377320: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1377320: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1377320: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1377320: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1377320: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1377320: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1377320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1377320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1377320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1380760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1380760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1380760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1382720: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1382720: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1382720: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1385000: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1385000: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1385000: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1385000: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1385000: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1385000: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1385000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1385000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1385000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1388440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1388440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1388440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1390400: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1390400: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1390400: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1392680: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1392680: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1392680: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1392680: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1392680: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1392680: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1392680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1392680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1392680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1396120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1396120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1396120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1398080: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1398080: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1398080: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1400360: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1400360: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1400360: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1400360: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1400360: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1400360: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1400360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1400360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1400360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1403800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1403800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1403800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1405760: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1405760: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1405760: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1408040: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1408040: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1408040: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1408040: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1408040: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1408040: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1408040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1408040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1408040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1411480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1411480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1411480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1413440: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1413440: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1413440: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1415720: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1415720: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1415720: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1415720: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1415720: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1415720: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1415720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1415720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1415720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1419160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1419160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1419160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1421120: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1421120: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1421120: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1423400: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1423400: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1423400: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1423400: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1423400: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1423400: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1423400: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1423400: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1423400: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1426840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1426840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1426840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1428800: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1428800: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1428800: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1431080: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1431080: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1431080: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1431080: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1431080: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1431080: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1431080: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1431080: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1431080: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1434520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1434520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1434520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1436480: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1436480: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1436480: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1438760: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1438760: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1438760: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1438760: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1438760: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1438760: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1438760: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1438760: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1438760: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1442200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1442200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1442200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1444160: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1444160: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1444160: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1446440: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1446440: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1446440: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1446440: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1446440: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1446440: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1446440: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1446440: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1446440: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1449880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1449880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1449880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1451840: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1451840: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1451840: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1454120: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1454120: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1454120: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1454120: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1454120: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1454120: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1454120: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1454120: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1454120: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1457560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1457560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1457560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1459520: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1459520: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1459520: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1461800: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1461800: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1461800: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1461800: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1461800: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1461800: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1461800: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1461800: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1461800: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1465240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1465240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1465240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1467200: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1467200: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1467200: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1469480: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1469480: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1469480: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1469480: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1469480: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1469480: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1469480: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1469480: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1469480: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1472920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1472920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1472920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1474880: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1474880: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1474880: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1477160: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1477160: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1477160: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1477160: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1477160: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1477160: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1477160: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1477160: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1477160: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1480600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1480600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1480600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1482560: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1482560: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1482560: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1484840: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1484840: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1484840: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1484840: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1484840: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1484840: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1484840: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1484840: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1484840: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1488280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1488280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1488280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1490240: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1490240: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1490240: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1492520: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1492520: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1492520: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1492520: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1492520: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1492520: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1492520: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1492520: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1492520: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1495960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1495960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1495960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1497920: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1497920: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1497920: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1500200: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1500200: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1500200: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1500200: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1500200: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1500200: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1500200: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1500200: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1500200: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1503640: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1503640: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1503640: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1505600: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1505600: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1505600: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1507880: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1507880: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1507880: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1507880: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1507880: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1507880: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1507880: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1507880: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1507880: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1511320: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1511320: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1511320: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1513280: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1513280: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1513280: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1515560: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1515560: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1515560: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1515560: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1515560: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1515560: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1515560: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1515560: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1515560: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1519000: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1519000: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1519000: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1520960: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1520960: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1520960: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1523240: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1523240: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1523240: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1523240: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1523240: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1523240: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1523240: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1523240: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1523240: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1526680: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1526680: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1526680: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1528640: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1528640: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1528640: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1530920: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1530920: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1530920: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1530920: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1530920: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1530920: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1530920: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1530920: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1530920: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1534360: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1534360: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1534360: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1536320: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1536320: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1536320: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1538600: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1538600: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1538600: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1538600: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1538600: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1538600: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1538600: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1538600: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1538600: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1542040: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1542040: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1542040: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1544000: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1544000: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1544000: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1546280: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1546280: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1546280: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1546280: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1546280: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1546280: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1546280: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1546280: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1546280: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(373) @ 1549720: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1549720: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1549720: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# UVM_INFO c_scoreboard.svh(251) @ 1551680: uvm_test_top.env.scoreboard [Report] transform y rightly
# UVM_INFO c_scoreboard.svh(256) @ 1551680: uvm_test_top.env.scoreboard [Report] transform cb rightly
# UVM_INFO c_scoreboard.svh(261) @ 1551680: uvm_test_top.env.scoreboard [Report] transform cr rightly
# UVM_INFO c_scoreboard.svh(304) @ 1553960: uvm_test_top.env.scoreboard [Report] fdct for y rightly
# UVM_INFO c_scoreboard.svh(310) @ 1553960: uvm_test_top.env.scoreboard [Report] fdct for cb rightly
# UVM_INFO c_scoreboard.svh(316) @ 1553960: uvm_test_top.env.scoreboard [Report] fdct for cr rightly
# UVM_INFO c_scoreboard.svh(278) @ 1553960: uvm_test_top.env.scoreboard [Report] quantize y rightly
# UVM_INFO c_scoreboard.svh(283) @ 1553960: uvm_test_top.env.scoreboard [Report] quantize cb rightly
# UVM_INFO c_scoreboard.svh(288) @ 1553960: uvm_test_top.env.scoreboard [Report] quantize cr rightly
# UVM_INFO c_scoreboard.svh(373) @ 1553960: uvm_test_top.env.scoreboard [Report] Right :), y component encoding
# UVM_INFO c_scoreboard.svh(353) @ 1553960: uvm_test_top.env.scoreboard [Report] Right :), cb component encoding
# UVM_INFO c_scoreboard.svh(332) @ 1553960: uvm_test_top.env.scoreboard [Report] Right :), cr component encoding
# Break key hit
# Simulation stop requested.
# Stopped at basic_modules.v line 51
# exit
# End time: 11:20:15 on Aug 29,2018, Elapsed time: 0:00:40
# Errors: 0, Warnings: 1
